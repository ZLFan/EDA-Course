module ceshi(sw17,ledr17);
input sw17;
output ledr17;
assign ledr17=sw17;
endmodule
