library verilog;
use verilog.vl_types.all;
entity spi_three_wire_test is
end spi_three_wire_test;
