rom_railgun_inst : rom_railgun PORT MAP (
		address	 => address_sig,
		inclock	 => inclock_sig,
		q	 => q_sig
	);
