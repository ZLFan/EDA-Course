module seven(clk,reset,row,col);
input clk;
input reset;
output reg [15:0] row; //��
output reg [3:0] col;//��
initial col=4'b0;
parameter [2:0]s1=000;
parameter [2:0]s2=001;
parameter [2:0]s3=010;
parameter [2:0]s4=011;
reg[6:0]data;
reg [2:0]current_state;
reg [2:0]next_state;

reg divi_50hz; 
reg [24:0] count_reg1; //����һ��25λ�ļ���ֵ
always@(posedge clk)
  if(count_reg1==25'd24999) //��50Mhz / 50hz��/ 2 - 1
    begin
      divi_50hz <= ~ divi_50hz; //�ߵ͵�ƽ��ת
      count_reg1 <= 25'd0; //����ֵ����
    end
  else
    begin 
      count_reg1 <= count_reg1 + 25'd1;
    end

always @(posedge clk)
begin
if (!reset) col<=4'b0;
 else 
 begin //���ü����������е� 16 �ֱ��룺0000-1111
 if(col<15) col<=col+1;
	     else col<=4'b0000;
end
end




//reg [2:0]count;
always@(posedge divi_50hz)
begin
 current_state<=next_state;
end

always@(posedge divi_50hz)
begin
 case(current_state)
  s1:next_state<=s2;
  s2:next_state<=s3;
  s3:next_state<=s4;
  s4:next_state<=s1;
  default:next_state<=s1;
 endcase
end

always@(posedge divi_50hz or negedge reset)
begin
 case(current_state)
  s1:
   begin 
    if (!reset) row<=16'b0;
	else
		begin
		case (col)
			4'b0000: row<=16'b0001000001000000; //�� 1 ��
			4'b0001: row<=16'b0001000010000000; //�� 2 ��
			4'b0010: row<=16'b0001000100000000; //3
			4'b0011: row<=16'b0001001111111111; //4
			4'b0100: row<=16'b0001110000000010; //5
			4'b0101: row<=16'b0011000010000010; //6
			4'b0110: row<=16'b1101000010000010; //7
			4'b0111: row<=16'b0001000010000010; //8
			4'b1000: row<=16'b0001000010000010; //9
			4'b1001: row<=16'b0001011111111110; //10
			4'b1010: row<=16'b0001000010000010; //11
			4'b1011: row<=16'b0001000010000010; //12
			4'b1100: row<=16'b0001000010000010; //13
			4'b1101: row<=16'b0001000010000010; //14
			4'b1110: row<=16'b0001000000000010; //15
			4'b1111: row<=16'b0000000000000000; //16
			default:row<=16'b0000000000000000;
		endcase
		end
   end
  s2:
   begin 
    if (!reset) row<=16'b0;
	else
		begin
		case (col)
			4'b0000: row<=16'b0000001000000000; //�� 1 ��
			4'b0001: row<=16'b0000001000000000; //�� 2 ��
			4'b0010: row<=16'b1000001000000000; //3
			4'b0011: row<=16'b1000001000000000; //4
			4'b0100: row<=16'b1000001000000000; //5
			4'b0101: row<=16'b1000001000000000; //6
			4'b0110: row<=16'b1000001000000000; //7
			4'b0111: row<=16'b1111111111111110; //8
			4'b1000: row<=16'b1000001000000000; //9
			4'b1001: row<=16'b1000001000000000; //10
			4'b1010: row<=16'b1000001000000000; //11
			4'b1011: row<=16'b1000001000000000; //12
			4'b1100: row<=16'b1000001000000000; //13
			4'b1101: row<=16'b0000001000000000; //14
			4'b1110: row<=16'b0000001000000000; //15
			4'b1111: row<=16'b0000000000000000; //16
			default:row<=16'b0000000000000000;
		endcase
		end
   end
  s3:
  begin 
    if (!reset) row<=16'b0;
	else
		begin
		case (col)
			4'b0000: row<=16'b0011111111110000; //�� 1 ��
			4'b0001: row<=16'b0010000000100000; //�� 2 ��
			4'b0010: row<=16'b0010000000100000; //3
			4'b0011: row<=16'b0011111111110010; //4
			4'b0100: row<=16'b0000000000001100; //5
			4'b0101: row<=16'b0011111111110000; //6
			4'b0110: row<=16'b0010001000010000; //7
			4'b0111: row<=16'b0010001001100000; //8
			4'b1000: row<=16'b0011111111111111; //9
			4'b1001: row<=16'b1010001010010000; //10
			4'b1010: row<=16'b0110001001100000; //11
			4'b1011: row<=16'b0011111111111111; //12
			4'b1100: row<=16'b0010001011000000; //13
			4'b1101: row<=16'b0010001000110000; //14
			4'b1110: row<=16'b0010000000010000; //15
			4'b1111: row<=16'b0000000000000000; //16
			default:row<=16'b0000000000000000;
		endcase
		end
   end
  s4:
   begin 
    if (!reset) row<=16'b0;
	else
		begin
		case (col)
			4'b0000: row<=16'b0000000000000000; //�� 1 ��
			4'b0001: row<=16'b0111111111100000; //�� 2 ��
			4'b0010: row<=16'b0100000001000000; //3
			4'b0011: row<=16'b0100000001000000; //4
			4'b0100: row<=16'b0111111111100000; //5
			4'b0101: row<=16'b0000000000001000; //6
			4'b0110: row<=16'b1000011000010000; //7
			4'b0111: row<=16'b1011101000100000; //8
			4'b1000: row<=16'b1000001001000000; //9
			4'b1001: row<=16'b1000001010000100; //10
			4'b1010: row<=16'b1000001100000010; //11
			4'b1011: row<=16'b1111111111111100; //12
			4'b1100: row<=16'b1000001000000000; //13
			4'b1101: row<=16'b1000001000000000; //14
			4'b1110: row<=16'b0000001000000000; //15
			4'b1111: row<=16'b0000000000000000; //16
			default:row<=16'b0000000000000000;
		endcase
		end
   end
  default:
  begin 
    if (!reset) row<=16'b0;
	else
		begin
		case (col)
			4'b0000: row<=16'b0010000000010000; //�� 1 ��
			4'b0001: row<=16'b0010000000010000; //�� 2 ��
			4'b0010: row<=16'b0010000000010000; //3
			4'b0011: row<=16'b0010001111010000; //4
			4'b0100: row<=16'b0010001001010000; //5
			4'b0101: row<=16'b1111101001010000; //6
			4'b0110: row<=16'b0010101001010000; //7
			4'b0111: row<=16'b0010111111111111; //8
			4'b1000: row<=16'b0010101001010000; //9
			4'b1001: row<=16'b1111101001010000; //10
			4'b1010: row<=16'b0010001001010000; //11
			4'b1011: row<=16'b0010001111010000; //12
			4'b1100: row<=16'b0010000000010000; //13
			4'b1101: row<=16'b0010000000010000; //14
			4'b1110: row<=16'b0101110001011000; //15
			4'b1111: row<=16'b0010000000010000; //16
			default:row<=16'b0000000000000000;
		endcase
		end
   end
 endcase
end
endmodule
