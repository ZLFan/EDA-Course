library verilog;
use verilog.vl_types.all;
entity divclk_vlg_tst is
end divclk_vlg_tst;
