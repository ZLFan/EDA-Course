module bigwork