library verilog;
use verilog.vl_types.all;
entity base1_vlg_tst is
end base1_vlg_tst;
