library verilog;
use verilog.vl_types.all;
entity spi_write_test is
end spi_write_test;
