module Keybord(clk,reset,clear,lockkey,pw0,pw1,pw2,pw3);
input clk;
input reset;
input clear;
input lockkey;
output [3:0]pw0;
output [3:0]pw1;
output [3:0]pw2;
output [3:0]pw3;
	
endmodule
