library verilog;
use verilog.vl_types.all;
entity I2C_write_test is
end I2C_write_test;
